VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wrapped_spell
  CLASS BLOCK ;
  FOREIGN wrapped_spell ;
  ORIGIN 0.000 0.000 ;
  SIZE 440.000 BY 440.000 ;
  PIN active
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 436.000 51.720 440.000 52.320 ;
    END
  END active
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 107.480 4.000 108.080 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 371.770 0.000 372.050 4.000 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 436.000 331.880 440.000 332.480 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 436.000 402.600 440.000 403.200 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.130 0.000 241.410 4.000 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.610 0.000 258.890 4.000 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.970 0.000 36.250 4.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 436.000 191.800 440.000 192.400 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 436.000 386.280 440.000 386.880 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.330 0.000 43.610 4.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.450 0.000 145.730 4.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.770 436.000 27.050 440.000 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.450 436.000 260.730 440.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 280.200 4.000 280.800 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 275.170 436.000 275.450 440.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 355.210 436.000 355.490 440.000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 382.200 4.000 382.800 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 399.370 436.000 399.650 440.000 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.890 436.000 60.170 440.000 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.290 0.000 262.570 4.000 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 436.000 429.800 440.000 430.400 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 436.000 272.040 440.000 272.640 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.810 0.000 245.090 4.000 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 393.080 4.000 393.680 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.040 4.000 102.640 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.370 0.000 123.650 4.000 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.530 436.000 282.810 440.000 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 274.760 4.000 275.360 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 436.000 99.320 440.000 99.920 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 340.040 4.000 340.640 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 362.570 436.000 362.850 440.000 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.970 0.000 197.250 4.000 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.250 436.000 136.530 440.000 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.570 436.000 293.850 440.000 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 297.250 436.000 297.530 440.000 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.410 436.000 88.690 440.000 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 419.610 0.000 419.890 4.000 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.530 436.000 52.810 440.000 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 335.890 0.000 336.170 4.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 436.000 29.960 440.000 30.560 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 178.200 4.000 178.800 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 436.000 277.480 440.000 278.080 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.970 436.000 312.250 440.000 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.850 436.000 49.130 440.000 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.090 436.000 184.370 440.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.090 0.000 299.370 4.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 436.000 342.760 440.000 343.360 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.170 436.000 114.450 440.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 365.880 4.000 366.480 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.810 436.000 38.090 440.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 426.970 0.000 427.250 4.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 178.570 0.000 178.850 4.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.250 436.000 67.530 440.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 390.170 0.000 390.450 4.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.210 436.000 56.490 440.000 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 140.120 4.000 140.720 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 334.600 4.000 335.200 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 436.000 104.760 440.000 105.360 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 258.440 4.000 259.040 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.090 0.000 230.370 4.000 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.010 436.000 392.290 440.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 436.000 115.640 440.000 116.240 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 350.610 0.000 350.890 4.000 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.210 436.000 286.490 440.000 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 376.760 4.000 377.360 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 278.850 436.000 279.130 440.000 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.160 4.000 193.760 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 436.000 391.720 440.000 392.320 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 436.000 129.170 440.000 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 379.130 0.000 379.410 4.000 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.130 436.000 34.410 440.000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.050 436.000 12.330 440.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 247.560 4.000 248.160 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 134.680 4.000 135.280 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.290 436.000 216.570 440.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 310.130 0.000 310.410 4.000 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 432.490 436.000 432.770 440.000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 436.000 282.920 440.000 283.520 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.690 436.000 73.970 440.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 304.610 436.000 304.890 440.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 371.320 4.000 371.920 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 436.600 4.000 437.200 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 436.000 418.920 440.000 419.520 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.850 436.000 118.130 440.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 256.770 436.000 257.050 440.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 15.000 4.000 15.600 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.770 0.000 73.050 4.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 403.960 4.000 404.560 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 436.000 180.920 440.000 181.520 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.920 4.000 113.520 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 58.520 4.000 59.120 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 397.530 0.000 397.810 4.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 291.080 4.000 291.680 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.970 0.000 358.250 4.000 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 436.000 375.400 440.000 376.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 436.000 68.040 440.000 68.640 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.210 0.000 171.490 4.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.050 436.000 81.330 440.000 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 253.090 436.000 253.370 440.000 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 436.000 293.800 440.000 294.400 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 340.490 436.000 340.770 440.000 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 345.480 4.000 346.080 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 343.250 0.000 343.530 4.000 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 130.730 0.000 131.010 4.000 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.010 436.000 162.290 440.000 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.690 436.000 234.970 440.000 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 421.450 436.000 421.730 440.000 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.890 436.000 198.170 440.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.010 436.000 70.290 440.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.930 436.000 140.210 440.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 253.000 4.000 253.600 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 436.000 2.760 440.000 3.360 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.090 436.000 92.370 440.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 415.930 0.000 416.210 4.000 ;
    END
  END io_out[9]
  PIN la1_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.490 436.000 271.770 440.000 ;
    END
  END la1_data_in[0]
  PIN la1_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.370 436.000 77.650 440.000 ;
    END
  END la1_data_in[10]
  PIN la1_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.330 436.000 158.610 440.000 ;
    END
  END la1_data_in[11]
  PIN la1_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.010 0.000 438.290 4.000 ;
    END
  END la1_data_in[12]
  PIN la1_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.370 0.000 215.650 4.000 ;
    END
  END la1_data_in[13]
  PIN la1_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 306.450 0.000 306.730 4.000 ;
    END
  END la1_data_in[14]
  PIN la1_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 436.000 24.520 440.000 25.120 ;
    END
  END la1_data_in[15]
  PIN la1_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 0.000 109.850 4.000 ;
    END
  END la1_data_in[16]
  PIN la1_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 434.330 0.000 434.610 4.000 ;
    END
  END la1_data_in[17]
  PIN la1_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 436.000 110.200 440.000 110.800 ;
    END
  END la1_data_in[18]
  PIN la1_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 384.650 436.000 384.930 440.000 ;
    END
  END la1_data_in[19]
  PIN la1_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 403.050 436.000 403.330 440.000 ;
    END
  END la1_data_in[1]
  PIN la1_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 436.000 408.040 440.000 408.640 ;
    END
  END la1_data_in[20]
  PIN la1_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 436.000 353.640 440.000 354.240 ;
    END
  END la1_data_in[21]
  PIN la1_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 332.210 0.000 332.490 4.000 ;
    END
  END la1_data_in[22]
  PIN la1_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.410 436.000 318.690 440.000 ;
    END
  END la1_data_in[23]
  PIN la1_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 167.320 4.000 167.920 ;
    END
  END la1_data_in[24]
  PIN la1_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.850 436.000 348.130 440.000 ;
    END
  END la1_data_in[25]
  PIN la1_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 373.610 436.000 373.890 440.000 ;
    END
  END la1_data_in[26]
  PIN la1_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 428.810 436.000 429.090 440.000 ;
    END
  END la1_data_in[27]
  PIN la1_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 436.000 435.240 440.000 435.840 ;
    END
  END la1_data_in[28]
  PIN la1_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.610 0.000 120.890 4.000 ;
    END
  END la1_data_in[29]
  PIN la1_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.530 0.000 167.810 4.000 ;
    END
  END la1_data_in[2]
  PIN la1_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 436.000 266.600 440.000 267.200 ;
    END
  END la1_data_in[30]
  PIN la1_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 318.280 4.000 318.880 ;
    END
  END la1_data_in[31]
  PIN la1_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 31.320 4.000 31.920 ;
    END
  END la1_data_in[3]
  PIN la1_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 333.130 436.000 333.410 440.000 ;
    END
  END la1_data_in[4]
  PIN la1_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.250 0.000 251.530 4.000 ;
    END
  END la1_data_in[5]
  PIN la1_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.050 0.000 219.330 4.000 ;
    END
  END la1_data_in[6]
  PIN la1_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.570 436.000 132.850 440.000 ;
    END
  END la1_data_in[7]
  PIN la1_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.650 0.000 269.930 4.000 ;
    END
  END la1_data_in[8]
  PIN la1_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.490 0.000 87.770 4.000 ;
    END
  END la1_data_in[9]
  PIN la1_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.010 436.000 231.290 440.000 ;
    END
  END la1_data_out[0]
  PIN la1_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.850 0.000 164.130 4.000 ;
    END
  END la1_data_out[10]
  PIN la1_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.720 4.000 86.320 ;
    END
  END la1_data_out[11]
  PIN la1_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 436.000 235.320 440.000 235.920 ;
    END
  END la1_data_out[12]
  PIN la1_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 436.000 19.080 440.000 19.680 ;
    END
  END la1_data_out[13]
  PIN la1_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 151.000 4.000 151.600 ;
    END
  END la1_data_out[14]
  PIN la1_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 237.450 0.000 237.730 4.000 ;
    END
  END la1_data_out[15]
  PIN la1_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.010 436.000 1.290 440.000 ;
    END
  END la1_data_out[16]
  PIN la1_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.050 0.000 127.330 4.000 ;
    END
  END la1_data_out[17]
  PIN la1_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.810 0.000 153.090 4.000 ;
    END
  END la1_data_out[18]
  PIN la1_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.730 0.000 62.010 4.000 ;
    END
  END la1_data_out[19]
  PIN la1_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 436.000 126.520 440.000 127.120 ;
    END
  END la1_data_out[1]
  PIN la1_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 231.240 4.000 231.840 ;
    END
  END la1_data_out[20]
  PIN la1_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.450 436.000 30.730 440.000 ;
    END
  END la1_data_out[21]
  PIN la1_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 225.800 4.000 226.400 ;
    END
  END la1_data_out[22]
  PIN la1_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.370 436.000 169.650 440.000 ;
    END
  END la1_data_out[23]
  PIN la1_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 436.000 45.450 440.000 ;
    END
  END la1_data_out[24]
  PIN la1_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 436.000 337.320 440.000 337.920 ;
    END
  END la1_data_out[25]
  PIN la1_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 414.090 436.000 414.370 440.000 ;
    END
  END la1_data_out[26]
  PIN la1_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 436.000 142.840 440.000 143.440 ;
    END
  END la1_data_out[27]
  PIN la1_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.890 436.000 290.170 440.000 ;
    END
  END la1_data_out[28]
  PIN la1_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 285.640 4.000 286.240 ;
    END
  END la1_data_out[29]
  PIN la1_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.250 0.000 113.530 4.000 ;
    END
  END la1_data_out[2]
  PIN la1_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 134.410 0.000 134.690 4.000 ;
    END
  END la1_data_out[30]
  PIN la1_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 436.000 93.880 440.000 94.480 ;
    END
  END la1_data_out[31]
  PIN la1_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 214.920 4.000 215.520 ;
    END
  END la1_data_out[3]
  PIN la1_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.650 436.000 154.930 440.000 ;
    END
  END la1_data_out[4]
  PIN la1_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.810 436.000 268.090 440.000 ;
    END
  END la1_data_out[5]
  PIN la1_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 436.000 310.120 440.000 310.720 ;
    END
  END la1_data_out[6]
  PIN la1_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 223.650 436.000 223.930 440.000 ;
    END
  END la1_data_out[7]
  PIN la1_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 436.000 369.960 440.000 370.560 ;
    END
  END la1_data_out[8]
  PIN la1_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 404.890 0.000 405.170 4.000 ;
    END
  END la1_data_out[9]
  PIN la1_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 377.290 436.000 377.570 440.000 ;
    END
  END la1_oenb[0]
  PIN la1_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 9.560 4.000 10.160 ;
    END
  END la1_oenb[10]
  PIN la1_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.890 0.000 106.170 4.000 ;
    END
  END la1_oenb[11]
  PIN la1_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 123.800 4.000 124.400 ;
    END
  END la1_oenb[12]
  PIN la1_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.290 0.000 193.570 4.000 ;
    END
  END la1_oenb[13]
  PIN la1_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.290 436.000 147.570 440.000 ;
    END
  END la1_oenb[14]
  PIN la1_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.690 0.000 50.970 4.000 ;
    END
  END la1_oenb[15]
  PIN la1_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.450 436.000 99.730 440.000 ;
    END
  END la1_oenb[16]
  PIN la1_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.490 0.000 156.770 4.000 ;
    END
  END la1_oenb[17]
  PIN la1_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.810 436.000 107.090 440.000 ;
    END
  END la1_oenb[18]
  PIN la1_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 425.720 4.000 426.320 ;
    END
  END la1_oenb[19]
  PIN la1_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.930 436.000 209.210 440.000 ;
    END
  END la1_oenb[1]
  PIN la1_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 420.280 4.000 420.880 ;
    END
  END la1_oenb[20]
  PIN la1_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 423.290 0.000 423.570 4.000 ;
    END
  END la1_oenb[21]
  PIN la1_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.890 0.000 175.170 4.000 ;
    END
  END la1_oenb[22]
  PIN la1_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.530 0.000 98.810 4.000 ;
    END
  END la1_oenb[23]
  PIN la1_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 436.000 304.680 440.000 305.280 ;
    END
  END la1_oenb[24]
  PIN la1_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 436.000 88.440 440.000 89.040 ;
    END
  END la1_oenb[25]
  PIN la1_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 365.330 0.000 365.610 4.000 ;
    END
  END la1_oenb[26]
  PIN la1_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.610 436.000 212.890 440.000 ;
    END
  END la1_oenb[27]
  PIN la1_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.170 436.000 344.450 440.000 ;
    END
  END la1_oenb[28]
  PIN la1_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.880 4.000 26.480 ;
    END
  END la1_oenb[29]
  PIN la1_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 387.640 4.000 388.240 ;
    END
  END la1_oenb[2]
  PIN la1_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.410 436.000 249.690 440.000 ;
    END
  END la1_oenb[30]
  PIN la1_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.250 0.000 21.530 4.000 ;
    END
  END la1_oenb[31]
  PIN la1_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.130 0.000 149.410 4.000 ;
    END
  END la1_oenb[3]
  PIN la1_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 36.760 4.000 37.360 ;
    END
  END la1_oenb[4]
  PIN la1_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.530 0.000 328.810 4.000 ;
    END
  END la1_oenb[5]
  PIN la1_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 398.520 4.000 399.120 ;
    END
  END la1_oenb[6]
  PIN la1_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.810 0.000 84.090 4.000 ;
    END
  END la1_oenb[7]
  PIN la1_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 324.850 0.000 325.130 4.000 ;
    END
  END la1_oenb[8]
  PIN la1_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 436.000 153.720 440.000 154.320 ;
    END
  END la1_oenb[9]
  PIN rambus_wb_ack_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.610 436.000 143.890 440.000 ;
    END
  END rambus_wb_ack_i
  PIN rambus_wb_adr_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 204.040 4.000 204.640 ;
    END
  END rambus_wb_adr_o[0]
  PIN rambus_wb_adr_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 242.120 4.000 242.720 ;
    END
  END rambus_wb_adr_o[1]
  PIN rambus_wb_adr_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.730 436.000 16.010 440.000 ;
    END
  END rambus_wb_adr_o[2]
  PIN rambus_wb_adr_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 176.730 436.000 177.010 440.000 ;
    END
  END rambus_wb_adr_o[3]
  PIN rambus_wb_adr_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.050 436.000 242.330 440.000 ;
    END
  END rambus_wb_adr_o[4]
  PIN rambus_wb_adr_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 436.000 8.200 440.000 8.800 ;
    END
  END rambus_wb_adr_o[5]
  PIN rambus_wb_adr_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 369.930 436.000 370.210 440.000 ;
    END
  END rambus_wb_adr_o[6]
  PIN rambus_wb_adr_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 436.000 251.640 440.000 252.240 ;
    END
  END rambus_wb_adr_o[7]
  PIN rambus_wb_adr_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 436.000 359.080 440.000 359.680 ;
    END
  END rambus_wb_adr_o[8]
  PIN rambus_wb_adr_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 198.600 4.000 199.200 ;
    END
  END rambus_wb_adr_o[9]
  PIN rambus_wb_clk_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.210 436.000 194.490 440.000 ;
    END
  END rambus_wb_clk_o
  PIN rambus_wb_cyc_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.850 0.000 95.130 4.000 ;
    END
  END rambus_wb_cyc_o
  PIN rambus_wb_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 313.810 0.000 314.090 4.000 ;
    END
  END rambus_wb_dat_i[0]
  PIN rambus_wb_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 209.480 4.000 210.080 ;
    END
  END rambus_wb_dat_i[10]
  PIN rambus_wb_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 436.000 35.400 440.000 36.000 ;
    END
  END rambus_wb_dat_i[11]
  PIN rambus_wb_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.930 436.000 439.210 440.000 ;
    END
  END rambus_wb_dat_i[12]
  PIN rambus_wb_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 226.410 0.000 226.690 4.000 ;
    END
  END rambus_wb_dat_i[13]
  PIN rambus_wb_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 436.000 137.400 440.000 138.000 ;
    END
  END rambus_wb_dat_i[14]
  PIN rambus_wb_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 436.000 83.000 440.000 83.600 ;
    END
  END rambus_wb_dat_i[15]
  PIN rambus_wb_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 436.000 261.160 440.000 261.760 ;
    END
  END rambus_wb_dat_i[16]
  PIN rambus_wb_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 436.000 186.360 440.000 186.960 ;
    END
  END rambus_wb_dat_i[17]
  PIN rambus_wb_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.330 436.000 227.610 440.000 ;
    END
  END rambus_wb_dat_i[18]
  PIN rambus_wb_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 436.000 197.240 440.000 197.840 ;
    END
  END rambus_wb_dat_i[19]
  PIN rambus_wb_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 4.000 21.040 ;
    END
  END rambus_wb_dat_i[1]
  PIN rambus_wb_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.490 0.000 317.770 4.000 ;
    END
  END rambus_wb_dat_i[20]
  PIN rambus_wb_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.370 0.000 54.650 4.000 ;
    END
  END rambus_wb_dat_i[21]
  PIN rambus_wb_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 350.920 4.000 351.520 ;
    END
  END rambus_wb_dat_i[22]
  PIN rambus_wb_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.050 0.000 288.330 4.000 ;
    END
  END rambus_wb_dat_i[23]
  PIN rambus_wb_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 393.850 0.000 394.130 4.000 ;
    END
  END rambus_wb_dat_i[24]
  PIN rambus_wb_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.210 436.000 125.490 440.000 ;
    END
  END rambus_wb_dat_i[25]
  PIN rambus_wb_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 307.400 4.000 308.000 ;
    END
  END rambus_wb_dat_i[26]
  PIN rambus_wb_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.370 436.000 238.650 440.000 ;
    END
  END rambus_wb_dat_i[27]
  PIN rambus_wb_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 414.840 4.000 415.440 ;
    END
  END rambus_wb_dat_i[28]
  PIN rambus_wb_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.210 0.000 102.490 4.000 ;
    END
  END rambus_wb_dat_i[29]
  PIN rambus_wb_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 436.000 213.560 440.000 214.160 ;
    END
  END rambus_wb_dat_i[2]
  PIN rambus_wb_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 321.170 0.000 321.450 4.000 ;
    END
  END rambus_wb_dat_i[30]
  PIN rambus_wb_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 161.880 4.000 162.480 ;
    END
  END rambus_wb_dat_i[31]
  PIN rambus_wb_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.410 0.000 65.690 4.000 ;
    END
  END rambus_wb_dat_i[3]
  PIN rambus_wb_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 436.000 170.040 440.000 170.640 ;
    END
  END rambus_wb_dat_i[4]
  PIN rambus_wb_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 187.720 4.000 188.320 ;
    END
  END rambus_wb_dat_i[5]
  PIN rambus_wb_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 436.000 424.360 440.000 424.960 ;
    END
  END rambus_wb_dat_i[6]
  PIN rambus_wb_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 436.000 348.200 440.000 348.800 ;
    END
  END rambus_wb_dat_i[7]
  PIN rambus_wb_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 436.000 326.440 440.000 327.040 ;
    END
  END rambus_wb_dat_i[8]
  PIN rambus_wb_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 436.000 321.000 440.000 321.600 ;
    END
  END rambus_wb_dat_i[9]
  PIN rambus_wb_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.930 0.000 186.210 4.000 ;
    END
  END rambus_wb_dat_o[0]
  PIN rambus_wb_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 410.410 436.000 410.690 440.000 ;
    END
  END rambus_wb_dat_o[10]
  PIN rambus_wb_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.210 0.000 10.490 4.000 ;
    END
  END rambus_wb_dat_o[11]
  PIN rambus_wb_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.850 0.000 3.130 4.000 ;
    END
  END rambus_wb_dat_o[12]
  PIN rambus_wb_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.730 436.000 85.010 440.000 ;
    END
  END rambus_wb_dat_o[13]
  PIN rambus_wb_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.610 0.000 189.890 4.000 ;
    END
  END rambus_wb_dat_o[14]
  PIN rambus_wb_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 375.450 0.000 375.730 4.000 ;
    END
  END rambus_wb_dat_o[15]
  PIN rambus_wb_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 436.170 436.000 436.450 440.000 ;
    END
  END rambus_wb_dat_o[16]
  PIN rambus_wb_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 408.570 0.000 408.850 4.000 ;
    END
  END rambus_wb_dat_o[17]
  PIN rambus_wb_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.970 436.000 220.250 440.000 ;
    END
  END rambus_wb_dat_o[18]
  PIN rambus_wb_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 356.360 4.000 356.960 ;
    END
  END rambus_wb_dat_o[19]
  PIN rambus_wb_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.090 0.000 69.370 4.000 ;
    END
  END rambus_wb_dat_o[1]
  PIN rambus_wb_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.170 0.000 160.450 4.000 ;
    END
  END rambus_wb_dat_o[20]
  PIN rambus_wb_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 388.330 436.000 388.610 440.000 ;
    END
  END rambus_wb_dat_o[21]
  PIN rambus_wb_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 145.560 4.000 146.160 ;
    END
  END rambus_wb_dat_o[22]
  PIN rambus_wb_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.090 0.000 138.370 4.000 ;
    END
  END rambus_wb_dat_o[23]
  PIN rambus_wb_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 409.400 4.000 410.000 ;
    END
  END rambus_wb_dat_o[24]
  PIN rambus_wb_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 436.000 148.280 440.000 148.880 ;
    END
  END rambus_wb_dat_o[25]
  PIN rambus_wb_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 436.000 246.200 440.000 246.800 ;
    END
  END rambus_wb_dat_o[26]
  PIN rambus_wb_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.690 0.000 280.970 4.000 ;
    END
  END rambus_wb_dat_o[27]
  PIN rambus_wb_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 80.280 4.000 80.880 ;
    END
  END rambus_wb_dat_o[28]
  PIN rambus_wb_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 361.650 0.000 361.930 4.000 ;
    END
  END rambus_wb_dat_o[29]
  PIN rambus_wb_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 436.000 229.880 440.000 230.480 ;
    END
  END rambus_wb_dat_o[2]
  PIN rambus_wb_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 329.450 436.000 329.730 440.000 ;
    END
  END rambus_wb_dat_o[30]
  PIN rambus_wb_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 4.120 4.000 4.720 ;
    END
  END rambus_wb_dat_o[31]
  PIN rambus_wb_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.010 0.000 277.290 4.000 ;
    END
  END rambus_wb_dat_o[3]
  PIN rambus_wb_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 406.730 436.000 407.010 440.000 ;
    END
  END rambus_wb_dat_o[4]
  PIN rambus_wb_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 401.210 0.000 401.490 4.000 ;
    END
  END rambus_wb_dat_o[5]
  PIN rambus_wb_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 300.930 436.000 301.210 440.000 ;
    END
  END rambus_wb_dat_o[6]
  PIN rambus_wb_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 339.570 0.000 339.850 4.000 ;
    END
  END rambus_wb_dat_o[7]
  PIN rambus_wb_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 323.720 4.000 324.320 ;
    END
  END rambus_wb_dat_o[8]
  PIN rambus_wb_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.010 0.000 47.290 4.000 ;
    END
  END rambus_wb_dat_o[9]
  PIN rambus_wb_rst_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 436.000 159.160 440.000 159.760 ;
    END
  END rambus_wb_rst_o
  PIN rambus_wb_sel_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.570 436.000 63.850 440.000 ;
    END
  END rambus_wb_sel_o[0]
  PIN rambus_wb_sel_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 436.000 240.760 440.000 241.360 ;
    END
  END rambus_wb_sel_o[1]
  PIN rambus_wb_sel_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.170 0.000 91.450 4.000 ;
    END
  END rambus_wb_sel_o[2]
  PIN rambus_wb_sel_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 346.930 0.000 347.210 4.000 ;
    END
  END rambus_wb_sel_o[3]
  PIN rambus_wb_stb_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 187.770 436.000 188.050 440.000 ;
    END
  END rambus_wb_stb_o
  PIN rambus_wb_we_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 395.690 436.000 395.970 440.000 ;
    END
  END rambus_wb_we_o
  PIN user_irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 53.080 4.000 53.680 ;
    END
  END user_irq[0]
  PIN user_irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.240 4.000 129.840 ;
    END
  END user_irq[1]
  PIN user_irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.250 436.000 205.530 440.000 ;
    END
  END user_irq[2]
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 427.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 427.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 427.280 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 427.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 427.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 427.280 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 430.650 0.000 430.930 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.970 436.000 151.250 440.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 436.000 77.560 440.000 78.160 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.090 436.000 322.370 440.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 245.730 436.000 246.010 440.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.130 436.000 103.410 440.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 0.000 32.570 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 204.330 0.000 204.610 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 436.000 288.360 440.000 288.960 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 436.000 257.080 440.000 257.680 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.770 0.000 234.050 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 312.840 4.000 313.440 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 436.000 62.600 440.000 63.200 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 354.290 0.000 354.570 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.200 4.000 42.800 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 301.960 4.000 302.560 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.010 0.000 208.290 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 295.410 0.000 295.690 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 436.000 13.640 440.000 14.240 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.530 436.000 121.810 440.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 96.600 4.000 97.200 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.650 0.000 39.930 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 201.570 436.000 201.850 440.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 436.000 208.120 440.000 208.720 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 436.000 413.480 440.000 414.080 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 63.960 4.000 64.560 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 220.360 4.000 220.960 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 436.000 121.080 440.000 121.680 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 284.370 0.000 284.650 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 358.890 436.000 359.170 440.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.330 0.000 273.610 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 269.320 4.000 269.920 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.570 0.000 17.850 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 369.010 0.000 369.290 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 436.000 40.840 440.000 41.440 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.450 436.000 191.730 440.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 436.000 364.520 440.000 365.120 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 431.160 4.000 431.760 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.410 436.000 19.690 440.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.370 436.000 8.650 440.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.890 0.000 14.170 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 69.400 4.000 70.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 436.000 175.480 440.000 176.080 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 211.690 0.000 211.970 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.160 4.000 91.760 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 417.770 436.000 418.050 440.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.770 436.000 96.050 440.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 236.680 4.000 237.280 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 436.000 219.000 440.000 219.600 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 425.130 436.000 425.410 440.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 329.160 4.000 329.760 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 436.000 73.480 440.000 74.080 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.930 0.000 255.210 4.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.970 436.000 381.250 440.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.690 436.000 165.970 440.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.930 0.000 117.210 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 436.000 224.440 440.000 225.040 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.770 0.000 303.050 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 436.000 57.160 440.000 57.760 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 296.520 4.000 297.120 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 382.810 0.000 383.090 4.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.250 0.000 182.530 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 436.000 131.960 440.000 132.560 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 366.250 436.000 366.530 440.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 436.000 380.840 440.000 381.440 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.490 0.000 386.770 4.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.610 0.000 28.890 4.000 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 436.000 202.680 440.000 203.280 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.530 0.000 6.810 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 436.000 397.160 440.000 397.760 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.530 436.000 351.810 440.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 412.250 0.000 412.530 4.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 336.810 436.000 337.090 440.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 156.440 4.000 157.040 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 172.760 4.000 173.360 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 247.570 0.000 247.850 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 291.730 0.000 292.010 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 263.880 4.000 264.480 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.090 436.000 23.370 440.000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.050 436.000 173.330 440.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 182.280 4.000 182.880 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.450 0.000 76.730 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.930 0.000 25.210 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.130 436.000 264.410 440.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.410 436.000 180.690 440.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.650 0.000 200.930 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.770 436.000 326.050 440.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 436.000 46.280 440.000 46.880 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 361.800 4.000 362.400 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 436.000 315.560 440.000 316.160 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.130 0.000 80.410 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.770 0.000 142.050 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 436.000 299.240 440.000 299.840 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.730 0.000 223.010 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.650 436.000 315.930 440.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 308.290 436.000 308.570 440.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.490 436.000 41.770 440.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.490 436.000 110.770 440.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.970 0.000 266.250 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 118.360 4.000 118.960 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.690 436.000 4.970 440.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 436.000 164.600 440.000 165.200 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 437.775 427.125 ;
      LAYER met1 ;
        RECT 0.070 5.140 439.230 427.280 ;
      LAYER met2 ;
        RECT 0.100 435.720 0.730 437.085 ;
        RECT 1.570 435.720 4.410 437.085 ;
        RECT 5.250 435.720 8.090 437.085 ;
        RECT 8.930 435.720 11.770 437.085 ;
        RECT 12.610 435.720 15.450 437.085 ;
        RECT 16.290 435.720 19.130 437.085 ;
        RECT 19.970 435.720 22.810 437.085 ;
        RECT 23.650 435.720 26.490 437.085 ;
        RECT 27.330 435.720 30.170 437.085 ;
        RECT 31.010 435.720 33.850 437.085 ;
        RECT 34.690 435.720 37.530 437.085 ;
        RECT 38.370 435.720 41.210 437.085 ;
        RECT 42.050 435.720 44.890 437.085 ;
        RECT 45.730 435.720 48.570 437.085 ;
        RECT 49.410 435.720 52.250 437.085 ;
        RECT 53.090 435.720 55.930 437.085 ;
        RECT 56.770 435.720 59.610 437.085 ;
        RECT 60.450 435.720 63.290 437.085 ;
        RECT 64.130 435.720 66.970 437.085 ;
        RECT 67.810 435.720 69.730 437.085 ;
        RECT 70.570 435.720 73.410 437.085 ;
        RECT 74.250 435.720 77.090 437.085 ;
        RECT 77.930 435.720 80.770 437.085 ;
        RECT 81.610 435.720 84.450 437.085 ;
        RECT 85.290 435.720 88.130 437.085 ;
        RECT 88.970 435.720 91.810 437.085 ;
        RECT 92.650 435.720 95.490 437.085 ;
        RECT 96.330 435.720 99.170 437.085 ;
        RECT 100.010 435.720 102.850 437.085 ;
        RECT 103.690 435.720 106.530 437.085 ;
        RECT 107.370 435.720 110.210 437.085 ;
        RECT 111.050 435.720 113.890 437.085 ;
        RECT 114.730 435.720 117.570 437.085 ;
        RECT 118.410 435.720 121.250 437.085 ;
        RECT 122.090 435.720 124.930 437.085 ;
        RECT 125.770 435.720 128.610 437.085 ;
        RECT 129.450 435.720 132.290 437.085 ;
        RECT 133.130 435.720 135.970 437.085 ;
        RECT 136.810 435.720 139.650 437.085 ;
        RECT 140.490 435.720 143.330 437.085 ;
        RECT 144.170 435.720 147.010 437.085 ;
        RECT 147.850 435.720 150.690 437.085 ;
        RECT 151.530 435.720 154.370 437.085 ;
        RECT 155.210 435.720 158.050 437.085 ;
        RECT 158.890 435.720 161.730 437.085 ;
        RECT 162.570 435.720 165.410 437.085 ;
        RECT 166.250 435.720 169.090 437.085 ;
        RECT 169.930 435.720 172.770 437.085 ;
        RECT 173.610 435.720 176.450 437.085 ;
        RECT 177.290 435.720 180.130 437.085 ;
        RECT 180.970 435.720 183.810 437.085 ;
        RECT 184.650 435.720 187.490 437.085 ;
        RECT 188.330 435.720 191.170 437.085 ;
        RECT 192.010 435.720 193.930 437.085 ;
        RECT 194.770 435.720 197.610 437.085 ;
        RECT 198.450 435.720 201.290 437.085 ;
        RECT 202.130 435.720 204.970 437.085 ;
        RECT 205.810 435.720 208.650 437.085 ;
        RECT 209.490 435.720 212.330 437.085 ;
        RECT 213.170 435.720 216.010 437.085 ;
        RECT 216.850 435.720 219.690 437.085 ;
        RECT 220.530 435.720 223.370 437.085 ;
        RECT 224.210 435.720 227.050 437.085 ;
        RECT 227.890 435.720 230.730 437.085 ;
        RECT 231.570 435.720 234.410 437.085 ;
        RECT 235.250 435.720 238.090 437.085 ;
        RECT 238.930 435.720 241.770 437.085 ;
        RECT 242.610 435.720 245.450 437.085 ;
        RECT 246.290 435.720 249.130 437.085 ;
        RECT 249.970 435.720 252.810 437.085 ;
        RECT 253.650 435.720 256.490 437.085 ;
        RECT 257.330 435.720 260.170 437.085 ;
        RECT 261.010 435.720 263.850 437.085 ;
        RECT 264.690 435.720 267.530 437.085 ;
        RECT 268.370 435.720 271.210 437.085 ;
        RECT 272.050 435.720 274.890 437.085 ;
        RECT 275.730 435.720 278.570 437.085 ;
        RECT 279.410 435.720 282.250 437.085 ;
        RECT 283.090 435.720 285.930 437.085 ;
        RECT 286.770 435.720 289.610 437.085 ;
        RECT 290.450 435.720 293.290 437.085 ;
        RECT 294.130 435.720 296.970 437.085 ;
        RECT 297.810 435.720 300.650 437.085 ;
        RECT 301.490 435.720 304.330 437.085 ;
        RECT 305.170 435.720 308.010 437.085 ;
        RECT 308.850 435.720 311.690 437.085 ;
        RECT 312.530 435.720 315.370 437.085 ;
        RECT 316.210 435.720 318.130 437.085 ;
        RECT 318.970 435.720 321.810 437.085 ;
        RECT 322.650 435.720 325.490 437.085 ;
        RECT 326.330 435.720 329.170 437.085 ;
        RECT 330.010 435.720 332.850 437.085 ;
        RECT 333.690 435.720 336.530 437.085 ;
        RECT 337.370 435.720 340.210 437.085 ;
        RECT 341.050 435.720 343.890 437.085 ;
        RECT 344.730 435.720 347.570 437.085 ;
        RECT 348.410 435.720 351.250 437.085 ;
        RECT 352.090 435.720 354.930 437.085 ;
        RECT 355.770 435.720 358.610 437.085 ;
        RECT 359.450 435.720 362.290 437.085 ;
        RECT 363.130 435.720 365.970 437.085 ;
        RECT 366.810 435.720 369.650 437.085 ;
        RECT 370.490 435.720 373.330 437.085 ;
        RECT 374.170 435.720 377.010 437.085 ;
        RECT 377.850 435.720 380.690 437.085 ;
        RECT 381.530 435.720 384.370 437.085 ;
        RECT 385.210 435.720 388.050 437.085 ;
        RECT 388.890 435.720 391.730 437.085 ;
        RECT 392.570 435.720 395.410 437.085 ;
        RECT 396.250 435.720 399.090 437.085 ;
        RECT 399.930 435.720 402.770 437.085 ;
        RECT 403.610 435.720 406.450 437.085 ;
        RECT 407.290 435.720 410.130 437.085 ;
        RECT 410.970 435.720 413.810 437.085 ;
        RECT 414.650 435.720 417.490 437.085 ;
        RECT 418.330 435.720 421.170 437.085 ;
        RECT 422.010 435.720 424.850 437.085 ;
        RECT 425.690 435.720 428.530 437.085 ;
        RECT 429.370 435.720 432.210 437.085 ;
        RECT 433.050 435.720 435.890 437.085 ;
        RECT 436.730 435.720 438.650 437.085 ;
        RECT 0.100 4.280 439.200 435.720 ;
        RECT 0.650 2.875 2.570 4.280 ;
        RECT 3.410 2.875 6.250 4.280 ;
        RECT 7.090 2.875 9.930 4.280 ;
        RECT 10.770 2.875 13.610 4.280 ;
        RECT 14.450 2.875 17.290 4.280 ;
        RECT 18.130 2.875 20.970 4.280 ;
        RECT 21.810 2.875 24.650 4.280 ;
        RECT 25.490 2.875 28.330 4.280 ;
        RECT 29.170 2.875 32.010 4.280 ;
        RECT 32.850 2.875 35.690 4.280 ;
        RECT 36.530 2.875 39.370 4.280 ;
        RECT 40.210 2.875 43.050 4.280 ;
        RECT 43.890 2.875 46.730 4.280 ;
        RECT 47.570 2.875 50.410 4.280 ;
        RECT 51.250 2.875 54.090 4.280 ;
        RECT 54.930 2.875 57.770 4.280 ;
        RECT 58.610 2.875 61.450 4.280 ;
        RECT 62.290 2.875 65.130 4.280 ;
        RECT 65.970 2.875 68.810 4.280 ;
        RECT 69.650 2.875 72.490 4.280 ;
        RECT 73.330 2.875 76.170 4.280 ;
        RECT 77.010 2.875 79.850 4.280 ;
        RECT 80.690 2.875 83.530 4.280 ;
        RECT 84.370 2.875 87.210 4.280 ;
        RECT 88.050 2.875 90.890 4.280 ;
        RECT 91.730 2.875 94.570 4.280 ;
        RECT 95.410 2.875 98.250 4.280 ;
        RECT 99.090 2.875 101.930 4.280 ;
        RECT 102.770 2.875 105.610 4.280 ;
        RECT 106.450 2.875 109.290 4.280 ;
        RECT 110.130 2.875 112.970 4.280 ;
        RECT 113.810 2.875 116.650 4.280 ;
        RECT 117.490 2.875 120.330 4.280 ;
        RECT 121.170 2.875 123.090 4.280 ;
        RECT 123.930 2.875 126.770 4.280 ;
        RECT 127.610 2.875 130.450 4.280 ;
        RECT 131.290 2.875 134.130 4.280 ;
        RECT 134.970 2.875 137.810 4.280 ;
        RECT 138.650 2.875 141.490 4.280 ;
        RECT 142.330 2.875 145.170 4.280 ;
        RECT 146.010 2.875 148.850 4.280 ;
        RECT 149.690 2.875 152.530 4.280 ;
        RECT 153.370 2.875 156.210 4.280 ;
        RECT 157.050 2.875 159.890 4.280 ;
        RECT 160.730 2.875 163.570 4.280 ;
        RECT 164.410 2.875 167.250 4.280 ;
        RECT 168.090 2.875 170.930 4.280 ;
        RECT 171.770 2.875 174.610 4.280 ;
        RECT 175.450 2.875 178.290 4.280 ;
        RECT 179.130 2.875 181.970 4.280 ;
        RECT 182.810 2.875 185.650 4.280 ;
        RECT 186.490 2.875 189.330 4.280 ;
        RECT 190.170 2.875 193.010 4.280 ;
        RECT 193.850 2.875 196.690 4.280 ;
        RECT 197.530 2.875 200.370 4.280 ;
        RECT 201.210 2.875 204.050 4.280 ;
        RECT 204.890 2.875 207.730 4.280 ;
        RECT 208.570 2.875 211.410 4.280 ;
        RECT 212.250 2.875 215.090 4.280 ;
        RECT 215.930 2.875 218.770 4.280 ;
        RECT 219.610 2.875 222.450 4.280 ;
        RECT 223.290 2.875 226.130 4.280 ;
        RECT 226.970 2.875 229.810 4.280 ;
        RECT 230.650 2.875 233.490 4.280 ;
        RECT 234.330 2.875 237.170 4.280 ;
        RECT 238.010 2.875 240.850 4.280 ;
        RECT 241.690 2.875 244.530 4.280 ;
        RECT 245.370 2.875 247.290 4.280 ;
        RECT 248.130 2.875 250.970 4.280 ;
        RECT 251.810 2.875 254.650 4.280 ;
        RECT 255.490 2.875 258.330 4.280 ;
        RECT 259.170 2.875 262.010 4.280 ;
        RECT 262.850 2.875 265.690 4.280 ;
        RECT 266.530 2.875 269.370 4.280 ;
        RECT 270.210 2.875 273.050 4.280 ;
        RECT 273.890 2.875 276.730 4.280 ;
        RECT 277.570 2.875 280.410 4.280 ;
        RECT 281.250 2.875 284.090 4.280 ;
        RECT 284.930 2.875 287.770 4.280 ;
        RECT 288.610 2.875 291.450 4.280 ;
        RECT 292.290 2.875 295.130 4.280 ;
        RECT 295.970 2.875 298.810 4.280 ;
        RECT 299.650 2.875 302.490 4.280 ;
        RECT 303.330 2.875 306.170 4.280 ;
        RECT 307.010 2.875 309.850 4.280 ;
        RECT 310.690 2.875 313.530 4.280 ;
        RECT 314.370 2.875 317.210 4.280 ;
        RECT 318.050 2.875 320.890 4.280 ;
        RECT 321.730 2.875 324.570 4.280 ;
        RECT 325.410 2.875 328.250 4.280 ;
        RECT 329.090 2.875 331.930 4.280 ;
        RECT 332.770 2.875 335.610 4.280 ;
        RECT 336.450 2.875 339.290 4.280 ;
        RECT 340.130 2.875 342.970 4.280 ;
        RECT 343.810 2.875 346.650 4.280 ;
        RECT 347.490 2.875 350.330 4.280 ;
        RECT 351.170 2.875 354.010 4.280 ;
        RECT 354.850 2.875 357.690 4.280 ;
        RECT 358.530 2.875 361.370 4.280 ;
        RECT 362.210 2.875 365.050 4.280 ;
        RECT 365.890 2.875 368.730 4.280 ;
        RECT 369.570 2.875 371.490 4.280 ;
        RECT 372.330 2.875 375.170 4.280 ;
        RECT 376.010 2.875 378.850 4.280 ;
        RECT 379.690 2.875 382.530 4.280 ;
        RECT 383.370 2.875 386.210 4.280 ;
        RECT 387.050 2.875 389.890 4.280 ;
        RECT 390.730 2.875 393.570 4.280 ;
        RECT 394.410 2.875 397.250 4.280 ;
        RECT 398.090 2.875 400.930 4.280 ;
        RECT 401.770 2.875 404.610 4.280 ;
        RECT 405.450 2.875 408.290 4.280 ;
        RECT 409.130 2.875 411.970 4.280 ;
        RECT 412.810 2.875 415.650 4.280 ;
        RECT 416.490 2.875 419.330 4.280 ;
        RECT 420.170 2.875 423.010 4.280 ;
        RECT 423.850 2.875 426.690 4.280 ;
        RECT 427.530 2.875 430.370 4.280 ;
        RECT 431.210 2.875 434.050 4.280 ;
        RECT 434.890 2.875 437.730 4.280 ;
        RECT 438.570 2.875 439.200 4.280 ;
      LAYER met3 ;
        RECT 4.400 436.240 436.000 437.065 ;
        RECT 4.400 436.200 435.600 436.240 ;
        RECT 4.000 434.840 435.600 436.200 ;
        RECT 4.000 432.160 436.000 434.840 ;
        RECT 4.400 430.800 436.000 432.160 ;
        RECT 4.400 430.760 435.600 430.800 ;
        RECT 4.000 429.400 435.600 430.760 ;
        RECT 4.000 426.720 436.000 429.400 ;
        RECT 4.400 425.360 436.000 426.720 ;
        RECT 4.400 425.320 435.600 425.360 ;
        RECT 4.000 423.960 435.600 425.320 ;
        RECT 4.000 421.280 436.000 423.960 ;
        RECT 4.400 419.920 436.000 421.280 ;
        RECT 4.400 419.880 435.600 419.920 ;
        RECT 4.000 418.520 435.600 419.880 ;
        RECT 4.000 415.840 436.000 418.520 ;
        RECT 4.400 414.480 436.000 415.840 ;
        RECT 4.400 414.440 435.600 414.480 ;
        RECT 4.000 413.080 435.600 414.440 ;
        RECT 4.000 410.400 436.000 413.080 ;
        RECT 4.400 409.040 436.000 410.400 ;
        RECT 4.400 409.000 435.600 409.040 ;
        RECT 4.000 407.640 435.600 409.000 ;
        RECT 4.000 404.960 436.000 407.640 ;
        RECT 4.400 403.600 436.000 404.960 ;
        RECT 4.400 403.560 435.600 403.600 ;
        RECT 4.000 402.200 435.600 403.560 ;
        RECT 4.000 399.520 436.000 402.200 ;
        RECT 4.400 398.160 436.000 399.520 ;
        RECT 4.400 398.120 435.600 398.160 ;
        RECT 4.000 396.760 435.600 398.120 ;
        RECT 4.000 394.080 436.000 396.760 ;
        RECT 4.400 392.720 436.000 394.080 ;
        RECT 4.400 392.680 435.600 392.720 ;
        RECT 4.000 391.320 435.600 392.680 ;
        RECT 4.000 388.640 436.000 391.320 ;
        RECT 4.400 387.280 436.000 388.640 ;
        RECT 4.400 387.240 435.600 387.280 ;
        RECT 4.000 385.880 435.600 387.240 ;
        RECT 4.000 383.200 436.000 385.880 ;
        RECT 4.400 381.840 436.000 383.200 ;
        RECT 4.400 381.800 435.600 381.840 ;
        RECT 4.000 380.440 435.600 381.800 ;
        RECT 4.000 377.760 436.000 380.440 ;
        RECT 4.400 376.400 436.000 377.760 ;
        RECT 4.400 376.360 435.600 376.400 ;
        RECT 4.000 375.000 435.600 376.360 ;
        RECT 4.000 372.320 436.000 375.000 ;
        RECT 4.400 370.960 436.000 372.320 ;
        RECT 4.400 370.920 435.600 370.960 ;
        RECT 4.000 369.560 435.600 370.920 ;
        RECT 4.000 366.880 436.000 369.560 ;
        RECT 4.400 365.520 436.000 366.880 ;
        RECT 4.400 365.480 435.600 365.520 ;
        RECT 4.000 364.120 435.600 365.480 ;
        RECT 4.000 362.800 436.000 364.120 ;
        RECT 4.400 361.400 436.000 362.800 ;
        RECT 4.000 360.080 436.000 361.400 ;
        RECT 4.000 358.680 435.600 360.080 ;
        RECT 4.000 357.360 436.000 358.680 ;
        RECT 4.400 355.960 436.000 357.360 ;
        RECT 4.000 354.640 436.000 355.960 ;
        RECT 4.000 353.240 435.600 354.640 ;
        RECT 4.000 351.920 436.000 353.240 ;
        RECT 4.400 350.520 436.000 351.920 ;
        RECT 4.000 349.200 436.000 350.520 ;
        RECT 4.000 347.800 435.600 349.200 ;
        RECT 4.000 346.480 436.000 347.800 ;
        RECT 4.400 345.080 436.000 346.480 ;
        RECT 4.000 343.760 436.000 345.080 ;
        RECT 4.000 342.360 435.600 343.760 ;
        RECT 4.000 341.040 436.000 342.360 ;
        RECT 4.400 339.640 436.000 341.040 ;
        RECT 4.000 338.320 436.000 339.640 ;
        RECT 4.000 336.920 435.600 338.320 ;
        RECT 4.000 335.600 436.000 336.920 ;
        RECT 4.400 334.200 436.000 335.600 ;
        RECT 4.000 332.880 436.000 334.200 ;
        RECT 4.000 331.480 435.600 332.880 ;
        RECT 4.000 330.160 436.000 331.480 ;
        RECT 4.400 328.760 436.000 330.160 ;
        RECT 4.000 327.440 436.000 328.760 ;
        RECT 4.000 326.040 435.600 327.440 ;
        RECT 4.000 324.720 436.000 326.040 ;
        RECT 4.400 323.320 436.000 324.720 ;
        RECT 4.000 322.000 436.000 323.320 ;
        RECT 4.000 320.600 435.600 322.000 ;
        RECT 4.000 319.280 436.000 320.600 ;
        RECT 4.400 317.880 436.000 319.280 ;
        RECT 4.000 316.560 436.000 317.880 ;
        RECT 4.000 315.160 435.600 316.560 ;
        RECT 4.000 313.840 436.000 315.160 ;
        RECT 4.400 312.440 436.000 313.840 ;
        RECT 4.000 311.120 436.000 312.440 ;
        RECT 4.000 309.720 435.600 311.120 ;
        RECT 4.000 308.400 436.000 309.720 ;
        RECT 4.400 307.000 436.000 308.400 ;
        RECT 4.000 305.680 436.000 307.000 ;
        RECT 4.000 304.280 435.600 305.680 ;
        RECT 4.000 302.960 436.000 304.280 ;
        RECT 4.400 301.560 436.000 302.960 ;
        RECT 4.000 300.240 436.000 301.560 ;
        RECT 4.000 298.840 435.600 300.240 ;
        RECT 4.000 297.520 436.000 298.840 ;
        RECT 4.400 296.120 436.000 297.520 ;
        RECT 4.000 294.800 436.000 296.120 ;
        RECT 4.000 293.400 435.600 294.800 ;
        RECT 4.000 292.080 436.000 293.400 ;
        RECT 4.400 290.680 436.000 292.080 ;
        RECT 4.000 289.360 436.000 290.680 ;
        RECT 4.000 287.960 435.600 289.360 ;
        RECT 4.000 286.640 436.000 287.960 ;
        RECT 4.400 285.240 436.000 286.640 ;
        RECT 4.000 283.920 436.000 285.240 ;
        RECT 4.000 282.520 435.600 283.920 ;
        RECT 4.000 281.200 436.000 282.520 ;
        RECT 4.400 279.800 436.000 281.200 ;
        RECT 4.000 278.480 436.000 279.800 ;
        RECT 4.000 277.080 435.600 278.480 ;
        RECT 4.000 275.760 436.000 277.080 ;
        RECT 4.400 274.360 436.000 275.760 ;
        RECT 4.000 273.040 436.000 274.360 ;
        RECT 4.000 271.640 435.600 273.040 ;
        RECT 4.000 270.320 436.000 271.640 ;
        RECT 4.400 268.920 436.000 270.320 ;
        RECT 4.000 267.600 436.000 268.920 ;
        RECT 4.000 266.200 435.600 267.600 ;
        RECT 4.000 264.880 436.000 266.200 ;
        RECT 4.400 263.480 436.000 264.880 ;
        RECT 4.000 262.160 436.000 263.480 ;
        RECT 4.000 260.760 435.600 262.160 ;
        RECT 4.000 259.440 436.000 260.760 ;
        RECT 4.400 258.080 436.000 259.440 ;
        RECT 4.400 258.040 435.600 258.080 ;
        RECT 4.000 256.680 435.600 258.040 ;
        RECT 4.000 254.000 436.000 256.680 ;
        RECT 4.400 252.640 436.000 254.000 ;
        RECT 4.400 252.600 435.600 252.640 ;
        RECT 4.000 251.240 435.600 252.600 ;
        RECT 4.000 248.560 436.000 251.240 ;
        RECT 4.400 247.200 436.000 248.560 ;
        RECT 4.400 247.160 435.600 247.200 ;
        RECT 4.000 245.800 435.600 247.160 ;
        RECT 4.000 243.120 436.000 245.800 ;
        RECT 4.400 241.760 436.000 243.120 ;
        RECT 4.400 241.720 435.600 241.760 ;
        RECT 4.000 240.360 435.600 241.720 ;
        RECT 4.000 237.680 436.000 240.360 ;
        RECT 4.400 236.320 436.000 237.680 ;
        RECT 4.400 236.280 435.600 236.320 ;
        RECT 4.000 234.920 435.600 236.280 ;
        RECT 4.000 232.240 436.000 234.920 ;
        RECT 4.400 230.880 436.000 232.240 ;
        RECT 4.400 230.840 435.600 230.880 ;
        RECT 4.000 229.480 435.600 230.840 ;
        RECT 4.000 226.800 436.000 229.480 ;
        RECT 4.400 225.440 436.000 226.800 ;
        RECT 4.400 225.400 435.600 225.440 ;
        RECT 4.000 224.040 435.600 225.400 ;
        RECT 4.000 221.360 436.000 224.040 ;
        RECT 4.400 220.000 436.000 221.360 ;
        RECT 4.400 219.960 435.600 220.000 ;
        RECT 4.000 218.600 435.600 219.960 ;
        RECT 4.000 215.920 436.000 218.600 ;
        RECT 4.400 214.560 436.000 215.920 ;
        RECT 4.400 214.520 435.600 214.560 ;
        RECT 4.000 213.160 435.600 214.520 ;
        RECT 4.000 210.480 436.000 213.160 ;
        RECT 4.400 209.120 436.000 210.480 ;
        RECT 4.400 209.080 435.600 209.120 ;
        RECT 4.000 207.720 435.600 209.080 ;
        RECT 4.000 205.040 436.000 207.720 ;
        RECT 4.400 203.680 436.000 205.040 ;
        RECT 4.400 203.640 435.600 203.680 ;
        RECT 4.000 202.280 435.600 203.640 ;
        RECT 4.000 199.600 436.000 202.280 ;
        RECT 4.400 198.240 436.000 199.600 ;
        RECT 4.400 198.200 435.600 198.240 ;
        RECT 4.000 196.840 435.600 198.200 ;
        RECT 4.000 194.160 436.000 196.840 ;
        RECT 4.400 192.800 436.000 194.160 ;
        RECT 4.400 192.760 435.600 192.800 ;
        RECT 4.000 191.400 435.600 192.760 ;
        RECT 4.000 188.720 436.000 191.400 ;
        RECT 4.400 187.360 436.000 188.720 ;
        RECT 4.400 187.320 435.600 187.360 ;
        RECT 4.000 185.960 435.600 187.320 ;
        RECT 4.000 183.280 436.000 185.960 ;
        RECT 4.400 181.920 436.000 183.280 ;
        RECT 4.400 181.880 435.600 181.920 ;
        RECT 4.000 180.520 435.600 181.880 ;
        RECT 4.000 179.200 436.000 180.520 ;
        RECT 4.400 177.800 436.000 179.200 ;
        RECT 4.000 176.480 436.000 177.800 ;
        RECT 4.000 175.080 435.600 176.480 ;
        RECT 4.000 173.760 436.000 175.080 ;
        RECT 4.400 172.360 436.000 173.760 ;
        RECT 4.000 171.040 436.000 172.360 ;
        RECT 4.000 169.640 435.600 171.040 ;
        RECT 4.000 168.320 436.000 169.640 ;
        RECT 4.400 166.920 436.000 168.320 ;
        RECT 4.000 165.600 436.000 166.920 ;
        RECT 4.000 164.200 435.600 165.600 ;
        RECT 4.000 162.880 436.000 164.200 ;
        RECT 4.400 161.480 436.000 162.880 ;
        RECT 4.000 160.160 436.000 161.480 ;
        RECT 4.000 158.760 435.600 160.160 ;
        RECT 4.000 157.440 436.000 158.760 ;
        RECT 4.400 156.040 436.000 157.440 ;
        RECT 4.000 154.720 436.000 156.040 ;
        RECT 4.000 153.320 435.600 154.720 ;
        RECT 4.000 152.000 436.000 153.320 ;
        RECT 4.400 150.600 436.000 152.000 ;
        RECT 4.000 149.280 436.000 150.600 ;
        RECT 4.000 147.880 435.600 149.280 ;
        RECT 4.000 146.560 436.000 147.880 ;
        RECT 4.400 145.160 436.000 146.560 ;
        RECT 4.000 143.840 436.000 145.160 ;
        RECT 4.000 142.440 435.600 143.840 ;
        RECT 4.000 141.120 436.000 142.440 ;
        RECT 4.400 139.720 436.000 141.120 ;
        RECT 4.000 138.400 436.000 139.720 ;
        RECT 4.000 137.000 435.600 138.400 ;
        RECT 4.000 135.680 436.000 137.000 ;
        RECT 4.400 134.280 436.000 135.680 ;
        RECT 4.000 132.960 436.000 134.280 ;
        RECT 4.000 131.560 435.600 132.960 ;
        RECT 4.000 130.240 436.000 131.560 ;
        RECT 4.400 128.840 436.000 130.240 ;
        RECT 4.000 127.520 436.000 128.840 ;
        RECT 4.000 126.120 435.600 127.520 ;
        RECT 4.000 124.800 436.000 126.120 ;
        RECT 4.400 123.400 436.000 124.800 ;
        RECT 4.000 122.080 436.000 123.400 ;
        RECT 4.000 120.680 435.600 122.080 ;
        RECT 4.000 119.360 436.000 120.680 ;
        RECT 4.400 117.960 436.000 119.360 ;
        RECT 4.000 116.640 436.000 117.960 ;
        RECT 4.000 115.240 435.600 116.640 ;
        RECT 4.000 113.920 436.000 115.240 ;
        RECT 4.400 112.520 436.000 113.920 ;
        RECT 4.000 111.200 436.000 112.520 ;
        RECT 4.000 109.800 435.600 111.200 ;
        RECT 4.000 108.480 436.000 109.800 ;
        RECT 4.400 107.080 436.000 108.480 ;
        RECT 4.000 105.760 436.000 107.080 ;
        RECT 4.000 104.360 435.600 105.760 ;
        RECT 4.000 103.040 436.000 104.360 ;
        RECT 4.400 101.640 436.000 103.040 ;
        RECT 4.000 100.320 436.000 101.640 ;
        RECT 4.000 98.920 435.600 100.320 ;
        RECT 4.000 97.600 436.000 98.920 ;
        RECT 4.400 96.200 436.000 97.600 ;
        RECT 4.000 94.880 436.000 96.200 ;
        RECT 4.000 93.480 435.600 94.880 ;
        RECT 4.000 92.160 436.000 93.480 ;
        RECT 4.400 90.760 436.000 92.160 ;
        RECT 4.000 89.440 436.000 90.760 ;
        RECT 4.000 88.040 435.600 89.440 ;
        RECT 4.000 86.720 436.000 88.040 ;
        RECT 4.400 85.320 436.000 86.720 ;
        RECT 4.000 84.000 436.000 85.320 ;
        RECT 4.000 82.600 435.600 84.000 ;
        RECT 4.000 81.280 436.000 82.600 ;
        RECT 4.400 79.880 436.000 81.280 ;
        RECT 4.000 78.560 436.000 79.880 ;
        RECT 4.000 77.160 435.600 78.560 ;
        RECT 4.000 75.840 436.000 77.160 ;
        RECT 4.400 74.480 436.000 75.840 ;
        RECT 4.400 74.440 435.600 74.480 ;
        RECT 4.000 73.080 435.600 74.440 ;
        RECT 4.000 70.400 436.000 73.080 ;
        RECT 4.400 69.040 436.000 70.400 ;
        RECT 4.400 69.000 435.600 69.040 ;
        RECT 4.000 67.640 435.600 69.000 ;
        RECT 4.000 64.960 436.000 67.640 ;
        RECT 4.400 63.600 436.000 64.960 ;
        RECT 4.400 63.560 435.600 63.600 ;
        RECT 4.000 62.200 435.600 63.560 ;
        RECT 4.000 59.520 436.000 62.200 ;
        RECT 4.400 58.160 436.000 59.520 ;
        RECT 4.400 58.120 435.600 58.160 ;
        RECT 4.000 56.760 435.600 58.120 ;
        RECT 4.000 54.080 436.000 56.760 ;
        RECT 4.400 52.720 436.000 54.080 ;
        RECT 4.400 52.680 435.600 52.720 ;
        RECT 4.000 51.320 435.600 52.680 ;
        RECT 4.000 48.640 436.000 51.320 ;
        RECT 4.400 47.280 436.000 48.640 ;
        RECT 4.400 47.240 435.600 47.280 ;
        RECT 4.000 45.880 435.600 47.240 ;
        RECT 4.000 43.200 436.000 45.880 ;
        RECT 4.400 41.840 436.000 43.200 ;
        RECT 4.400 41.800 435.600 41.840 ;
        RECT 4.000 40.440 435.600 41.800 ;
        RECT 4.000 37.760 436.000 40.440 ;
        RECT 4.400 36.400 436.000 37.760 ;
        RECT 4.400 36.360 435.600 36.400 ;
        RECT 4.000 35.000 435.600 36.360 ;
        RECT 4.000 32.320 436.000 35.000 ;
        RECT 4.400 30.960 436.000 32.320 ;
        RECT 4.400 30.920 435.600 30.960 ;
        RECT 4.000 29.560 435.600 30.920 ;
        RECT 4.000 26.880 436.000 29.560 ;
        RECT 4.400 25.520 436.000 26.880 ;
        RECT 4.400 25.480 435.600 25.520 ;
        RECT 4.000 24.120 435.600 25.480 ;
        RECT 4.000 21.440 436.000 24.120 ;
        RECT 4.400 20.080 436.000 21.440 ;
        RECT 4.400 20.040 435.600 20.080 ;
        RECT 4.000 18.680 435.600 20.040 ;
        RECT 4.000 16.000 436.000 18.680 ;
        RECT 4.400 14.640 436.000 16.000 ;
        RECT 4.400 14.600 435.600 14.640 ;
        RECT 4.000 13.240 435.600 14.600 ;
        RECT 4.000 10.560 436.000 13.240 ;
        RECT 4.400 9.200 436.000 10.560 ;
        RECT 4.400 9.160 435.600 9.200 ;
        RECT 4.000 7.800 435.600 9.160 ;
        RECT 4.000 5.120 436.000 7.800 ;
        RECT 4.400 3.760 436.000 5.120 ;
        RECT 4.400 3.720 435.600 3.760 ;
        RECT 4.000 2.895 435.600 3.720 ;
      LAYER met4 ;
        RECT 76.655 10.240 97.440 376.545 ;
        RECT 99.840 10.240 174.240 376.545 ;
        RECT 176.640 10.240 251.040 376.545 ;
        RECT 253.440 10.240 327.840 376.545 ;
        RECT 330.240 10.240 404.640 376.545 ;
        RECT 407.040 10.240 421.985 376.545 ;
        RECT 76.655 8.335 421.985 10.240 ;
  END
END wrapped_spell
END LIBRARY

